//03/23/21 13:58:58
//Author��xuhao Yang
module  my_test();
    input 
    output

endmodule
